// File: matrix_multiply.v
module matrix_multiply (
    input clk,
    input rst,
    input start,
    input [31:0] A [0:3][0:3],
    input [31:0] B [0:3][0:3],
    output reg [31:0] C [0:3][0:3],
    output reg done
);

// RTL code for matrix multiplication which i really dont know 

endmodule
